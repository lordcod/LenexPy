<?xml version="1.0" encoding="utf-8"?>
<LENEX version="3.0">
    <CONSTRUCTOR name="Name" registration="Sport-Sbor Agency" version="11.80519">
        <CONTACT city="Spiegel b. Bern" country="CH" email="sales@swimrankings.net"
            internet="https://www.swimrankings.net" name="Splash Software GmbH" street="Ahornweg 41"
            zip="3095" />
    </CONSTRUCTOR>
    <MEETS>
        <MEET city="Наро-Фоминск" course="SCM" name="Свим Драйв " nation="RUS" timing="MANUAL1">
            <AGEDATE type="YEAR" value="2025-02-02" />
            <CLUBS>
                <CLUB name="Обнинск" nation="RUS" type="CLUB">
                    <CONTACT name="Обнинск" />
                    <ATHLETES>
                        <ATHLETE athleteid="1569" birthdate="2013-10-21" firstname="Даниил"
                            gender="M" lastname="Зыболов" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:16.00" eventid="1093" heatid="1809" lane="2" />
                                <ENTRY entrytime="00:00:17.00" eventid="1099" heatid="1813" lane="2" />
                                <ENTRY entrytime="00:00:34.00" eventid="1112" heatid="1829" lane="2" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1550" birthdate="2014-08-20" firstname="Назар"
                            gender="M" lastname="Киселев" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:19.00" eventid="1099" heatid="1813" lane="3" />
                                <ENTRY entrytime="00:00:35.00" eventid="1103" heatid="1822" lane="1" />
                                <ENTRY entrytime="00:00:38.00" eventid="1112" heatid="1829" lane="3" />
                            </ENTRIES>
                        </ATHLETE>
                    </ATHLETES>
                </CLUB>
                <CLUB name="Клин" nation="RUS" type="CLUB">
                    <CONTACT name="Клин" />
                    <ATHLETES>
                        <ATHLETE athleteid="1493" birthdate="2016-04-26" firstname="Злата"
                            gender="F" lastname="Крятова" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:34.50" eventid="1095" heatid="1810" lane="2" />
                                <ENTRY entrytime="00:00:47.40" eventid="1101" heatid="1815" lane="3" />
                                <ENTRY entrytime="00:00:33.30" eventid="1087" heatid="1803" lane="3" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1482" birthdate="2014-07-09" firstname="Изабелла"
                            gender="F" lastname="Крятова" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:43.00" eventid="1114" heatid="1830" lane="2" />
                                <ENTRY entrytime="00:00:23.00" eventid="1095" heatid="1811" lane="1" />
                                <ENTRY entrytime="00:00:40.00" eventid="1101" heatid="1816" lane="1" />
                            </ENTRIES>
                        </ATHLETE>
                    </ATHLETES>
                </CLUB>
                <CLUB name="Подольск" nation="RUS" type="CLUB">
                    <CONTACT name="Подольск" />
                    <ATHLETES>
                        <ATHLETE athleteid="1565" birthdate="2015-03-04" firstname="Алиса"
                            gender="F" lastname="Усманова" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="NT" eventid="1101" heatid="1814" lane="1" />
                                <ENTRY entrytime="NT" eventid="1110" heatid="1826" lane="4" />
                                <ENTRY entrytime="NT" eventid="1114" heatid="1830" lane="1" />
                            </ENTRIES>
                        </ATHLETE>
                    </ATHLETES>
                </CLUB>
                <CLUB name="ДЮСШ &quot;Воробьевы горы&quot;" nation="RUS" type="CLUB">
                    <ATHLETES>
                        <ATHLETE athleteid="1678" birthdate="2014-03-26" firstname="Ольга"
                            gender="F" lastname="Поздяева" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="NT" eventid="1087" heatid="1802" lane="2" />
                                <ENTRY entrytime="NT" eventid="1091" heatid="1805" lane="3" />
                                <ENTRY entrytime="NT" eventid="1095" heatid="1810" lane="3" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1683" birthdate="2014-03-26" firstname="Анастасия"
                            gender="F" lastname="Поздяева" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="NT" eventid="1087" heatid="1802" lane="3" />
                                <ENTRY entrytime="NT" eventid="1091" heatid="1805" lane="1" />
                                <ENTRY entrytime="NT" eventid="1095" heatid="1810" lane="1" />
                            </ENTRIES>
                        </ATHLETE>
                    </ATHLETES>
                </CLUB>
                <CLUB name="Фрязино" nation="RUS" type="CLUB">
                    <CONTACT name="Фрязино" />
                    <ATHLETES>
                        <ATHLETE athleteid="1585" birthdate="2019-01-15" firstname="Елизавета"
                            gender="F" lastname="Шкурак" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:01:47.09" eventid="1110" heatid="1826" lane="1" />
                                <ENTRY entrytime="00:00:53.04" eventid="1091" heatid="1805" lane="2" />
                                <ENTRY entrytime="00:00:48.05" eventid="1074" heatid="1800" lane="2" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1581" birthdate="2013-02-21" firstname="Матвей"
                            gender="M" lastname="Шкурак" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:22.05" eventid="1093" heatid="1809" lane="3" />
                                <ENTRY entrytime="00:00:38.09" eventid="1103" heatid="1821" lane="2" />
                                <ENTRY entrytime="00:00:25.03" eventid="1099" heatid="1813" lane="1" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1507" birthdate="2013-07-16" firstname="Ксения"
                            gender="F" lastname="Щербакова" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:17.00" eventid="1095" heatid="1811" lane="2" />
                                <ENTRY entrytime="00:00:45.00" eventid="1105" heatid="1823" lane="2" />
                                <ENTRY entrytime="00:00:43.00" eventid="1114" heatid="1830" lane="3" />
                            </ENTRIES>
                        </ATHLETE>
                    </ATHLETES>
                </CLUB>
                <CLUB name="Наро-Фоминск" nation="RUS" type="CLUB">
                    <CONTACT name="Наро-Фоминск" />
                    <ATHLETES>
                        <ATHLETE athleteid="1479" birthdate="2014-08-11" firstname="Захар"
                            gender="M" lastname="Бабичев" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:34.12" eventid="1103" heatid="1822" lane="3" />
                                <ENTRY entrytime="00:00:50.33" eventid="1107" heatid="1825" lane="3" />
                                <ENTRY entrytime="00:00:43.32" eventid="1116" heatid="1831" lane="2" />
                                <ENTRY entrytime="NT" eventid="1133" heatid="1833" lane="3">
                                    <MEETINFO qualificationtime="00:00:00.00" />
                                </ENTRY>
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1541" birthdate="2014-02-08" firstname="Ева" gender="F"
                            lastname="Хорошилова" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:01:30.00" eventid="1101" heatid="1814" lane="3"
                                    status="DNS" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1526" birthdate="2014-09-16" firstname="Иван" gender="M"
                            lastname="Губанов" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="NT" eventid="1103" heatid="1817" lane="2" />
                                <ENTRY entrytime="NT" eventid="1112" heatid="1827" lane="1" />
                                <ENTRY entrytime="NT" eventid="1107" heatid="1824" lane="3" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1515" birthdate="2013-05-17" firstname="Кирилл"
                            gender="M" lastname="Сердюков" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="NT" eventid="1103" heatid="1818" lane="2" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1561" birthdate="2015-12-17" firstname="Ярослав"
                            gender="M" lastname="Осипцов" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:01:00.00" eventid="1103" heatid="1819" lane="2" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1487" birthdate="2015-05-30" firstname="Захар"
                            gender="M" lastname="Рыбкин" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:45.53" eventid="1103" heatid="1821" lane="3" />
                                <ENTRY entrytime="00:00:50.23" eventid="1112" heatid="1829" lane="4" />
                                <ENTRY entrytime="NT" eventid="1089" heatid="1804" lane="1" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1549" birthdate="2012-07-23" firstname="Артём"
                            gender="M" lastname="Терёшкин" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:34.00" eventid="1103" heatid="1822" lane="2" />
                                <ENTRY entrytime="00:00:45.00" eventid="1107" heatid="1825" lane="2" />
                                <ENTRY entrytime="00:00:40.35" eventid="1112" heatid="1829" lane="1" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1555" birthdate="2007-05-12" firstname="Фёдор"
                            gender="M" lastname="Шарканов" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="NT" eventid="1121" heatid="1832" lane="3" />
                                <ENTRY entrytime="NT" eventid="1133" heatid="1833" lane="1">
                                    <MEETINFO qualificationtime="00:00:00.00" />
                                </ENTRY>
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1531" birthdate="2011-11-03" firstname="Леонид"
                            gender="M" lastname="Емельянов" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="NT" eventid="1093" heatid="1807" lane="1" />
                                <ENTRY entrytime="NT" eventid="1103" heatid="1818" lane="3" />
                                <ENTRY entrytime="NT" eventid="1099" heatid="1812" lane="3" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1574" birthdate="2016-07-12" firstname="Иван" gender="M"
                            lastname="Ишин" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:01:00.00" eventid="1085" heatid="1801" lane="2" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1529" birthdate="2014-12-28" firstname="Александр"
                            gender="M" lastname="Емельянов" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="NT" eventid="1103" heatid="1818" lane="1" />
                                <ENTRY entrytime="NT" eventid="1089" heatid="1804" lane="4" />
                                <ENTRY entrytime="NT" eventid="1093" heatid="1807" lane="2" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1671" birthdate="2017-03-24" firstname="Мирон"
                            gender="M" lastname="Шарканов" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="NT" eventid="1093" heatid="1807" lane="3" />
                                <ENTRY entrytime="NT" eventid="1112" heatid="1827" lane="3" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1552" birthdate="2012-03-05" firstname="Семён"
                            gender="M" lastname="Гришаев" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:47.00" eventid="1103" heatid="1821" lane="1" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1579" birthdate="2010-08-29" firstname="Евгений"
                            gender="M" lastname="Аверьянов" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:01:00.00" eventid="1103" heatid="1819" lane="3"
                                    status="DNS" />
                                <ENTRY entrytime="00:01:00.00" eventid="1112" heatid="1828" lane="1"
                                    status="DNS" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1519" birthdate="2019-03-26" firstname="Ярослав"
                            gender="M" lastname="Шавергин" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="NT" eventid="1085" heatid="1801" lane="3" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1798" birthdate="2016-08-03" firstname="Михаил"
                            gender="M" lastname="Шубин" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:50.00" eventid="1103" heatid="1821" lane="4" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1560" birthdate="2013-03-27" firstname="Вадим"
                            gender="M" lastname="Пушкарев" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:01:00.00" eventid="1103" heatid="1820" lane="4" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1491" birthdate="2010-08-11" firstname="Екатерина"
                            gender="F" lastname="Белых" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:32.20" eventid="1101" heatid="1816" lane="3" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1533" birthdate="2015-01-14" firstname="Марк" gender="M"
                            lastname="Фильчугов" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:58.09" eventid="1103" heatid="1820" lane="1" />
                                <ENTRY entrytime="00:00:59.08" eventid="1107" heatid="1825" lane="1" />
                                <ENTRY entrytime="00:00:59.09" eventid="1112" heatid="1828" lane="3" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1545" birthdate="2014-11-15" firstname="Владислав"
                            gender="M" lastname="Полуботко" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="NT" eventid="1103" heatid="1817" lane="1" />
                                <ENTRY entrytime="NT" eventid="1107" heatid="1824" lane="1" />
                                <ENTRY entrytime="NT" eventid="1112" heatid="1827" lane="2" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1477" birthdate="2014-01-27" firstname="Матвей"
                            gender="M" lastname="Скворцов" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:55.00" eventid="1103" heatid="1820" lane="3"
                                    status="DNS" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1556" birthdate="2016-08-23" firstname="Кирилл"
                            gender="M" lastname="Паспортников" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="NT" eventid="1103" heatid="1817" lane="3" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1535" birthdate="2014-08-10" firstname="Эмиль"
                            gender="M" lastname="Рожков" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:58.03" eventid="1089" heatid="1804" lane="3" />
                                <ENTRY entrytime="00:01:00.06" eventid="1107" heatid="1824" lane="2" />
                                <ENTRY entrytime="00:00:58.07" eventid="1093" heatid="1808" lane="1" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1497" birthdate="2016-08-04" firstname="Вероника"
                            gender="F" lastname="Жмуренко" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:01:30.00" eventid="1101" heatid="1814" lane="2" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1539" birthdate="2014-10-04" firstname="Андрей"
                            gender="M" lastname="Шишмарев" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:35.06" eventid="1103" heatid="1822" lane="4" />
                                <ENTRY entrytime="00:00:30.02" eventid="1093" heatid="1808" lane="2" />
                                <ENTRY entrytime="00:00:31.02" eventid="1089" heatid="1804" lane="2" />
                            </ENTRIES>
                        </ATHLETE>
                    </ATHLETES>
                </CLUB>
                <CLUB name="Москва" nation="RUS" type="CLUB">
                    <CONTACT name="Москва" />
                    <ATHLETES>
                        <ATHLETE athleteid="1505" birthdate="1975-03-20" firstname="Денис"
                            gender="M" lastname="Фокин" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="NT" eventid="1121" heatid="1832" lane="2" />
                                <ENTRY entrytime="NT" eventid="1133" heatid="1833" lane="2" />
                            </ENTRIES>
                        </ATHLETE>
                        <ATHLETE athleteid="1523" birthdate="2014-07-10" firstname="Андрей"
                            gender="M" lastname="Трофимов" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:53.73" eventid="1103" heatid="1820" lane="2" />
                                <ENTRY entrytime="NT" eventid="1099" heatid="1812" lane="2" />
                            </ENTRIES>
                        </ATHLETE>
                    </ATHLETES>
                </CLUB>
                <CLUB name="Дубна" nation="RUS" type="CLUB">
                    <CONTACT name="Дубна" />
                    <ATHLETES>
                        <ATHLETE athleteid="1516" birthdate="2017-06-26" firstname="Таисия"
                            gender="F" lastname="Большова" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:49.00" eventid="1101" heatid="1815" lane="1" />
                                <ENTRY entrytime="00:00:27.00" eventid="1087" heatid="1803" lane="2" />
                                <ENTRY entrytime="00:00:48.00" eventid="1110" heatid="1826" lane="2" />
                            </ENTRIES>
                        </ATHLETE>
                    </ATHLETES>
                </CLUB>
                <CLUB name="Бронницы" nation="RUS" type="CLUB">
                    <CONTACT name="Бронницы" />
                    <ATHLETES>
                        <ATHLETE athleteid="1674" birthdate="2017-06-06" firstname="Игорь"
                            gender="M" lastname="Орлов" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:23.00" eventid="1093" heatid="1809" lane="1" />
                                <ENTRY entrytime="00:00:56.00" eventid="1112" heatid="1828" lane="2" />
                                <ENTRY entrytime="00:01:45.00" eventid="1103" heatid="1819" lane="4" />
                            </ENTRIES>
                        </ATHLETE>
                    </ATHLETES>
                </CLUB>
                <CLUB name="Мытищи" nation="RUS" type="CLUB">
                    <CONTACT name="Мытищи" />
                    <ATHLETES>
                        <ATHLETE athleteid="1503" birthdate="2018-02-23" firstname="Артем"
                            gender="M" lastname="Литвинов" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:01:01.00" eventid="1103" heatid="1819" lane="1" />
                                <ENTRY entrytime="00:01:01.47" eventid="1112" heatid="1828" lane="4" />
                                <ENTRY entrytime="00:00:34.31" eventid="1093" heatid="1808" lane="3" />
                            </ENTRIES>
                        </ATHLETE>
                    </ATHLETES>
                </CLUB>
                <CLUB name="Воскресенск" nation="RUS" type="CLUB">
                    <CONTACT name="Воскресенск" />
                    <ATHLETES>
                        <ATHLETE athleteid="1502" birthdate="2019-05-12" firstname="Варвара"
                            gender="F" lastname="Шарина" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:45.00" eventid="1087" heatid="1803" lane="1" />
                                <ENTRY entrytime="00:00:35.00" eventid="1091" heatid="1806" lane="1" />
                            </ENTRIES>
                        </ATHLETE>
                    </ATHLETES>
                </CLUB>
                <CLUB name="Молодежный" nation="RUS" type="CLUB">
                    <CONTACT name="Молодежный" />
                    <ATHLETES>
                        <ATHLETE athleteid="1589" birthdate="2011-12-28" firstname="Олеся"
                            gender="F" lastname="Шевченко" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:19.30" eventid="1091" heatid="1806" lane="3" />
                                <ENTRY entrytime="00:00:32.11" eventid="1101" heatid="1816" lane="2" />
                                <ENTRY entrytime="00:00:19.30" eventid="1095" heatid="1811" lane="3" />
                            </ENTRIES>
                        </ATHLETE>
                    </ATHLETES>
                </CLUB>
                <CLUB name="Химки" nation="RUS" type="CLUB">
                    <CONTACT name="Химки" />
                    <ATHLETES>
                        <ATHLETE athleteid="1509" birthdate="2015-01-09" firstname="Ева" gender="F"
                            lastname="Горшкова" nation="RUS">
                            <ENTRIES>
                                <ENTRY entrytime="00:00:43.50" eventid="1101" heatid="1815" lane="2" />
                                <ENTRY entrytime="00:00:19.20" eventid="1091" heatid="1806" lane="2" />
                                <ENTRY entrytime="00:00:48.50" eventid="1110" heatid="1826" lane="3" />
                            </ENTRIES>
                        </ATHLETE>
                    </ATHLETES>
                </CLUB>
            </CLUBS>
            <POINTTABLE name="AQUA Point Scoring" pointtableid="3017" version="2024" />
            <POOL lanemax="4" lanemin="1" />
            <SESSIONS>
                <SESSION date="2025-02-02T00:00:00" daytime="10:30:00" number="1"
                    warmupfrom="10:00:00">
                    <EVENTS>
                        <EVENT daytime="10:30:00" eventid="1074" gender="F" number="1" order="1"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1075" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1135" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1136" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1137" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1138" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1139" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1140" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1141" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1142" agemax="14" agemin="14" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="10:30:00" heatid="1800" number="1" order="1"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE code="25 с дс" distance="25" name="25m На груди с доской"
                                relaycount="1" stroke="UNKNOWN" swimstyleid="101" />
                        </EVENT>
                        <EVENT daytime="10:30:00" eventid="1085" gender="M" number="2" order="2"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1143" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1144" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1145" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1146" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1147" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1148" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1149" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1150" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1151" agemax="14" agemin="14" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="10:30:00" heatid="1801" number="1" order="1"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE code="25 с дс" distance="25" name="25m На груди с доской"
                                relaycount="1" stroke="UNKNOWN" swimstyleid="101" />
                        </EVENT>
                        <EVENT daytime="10:35:00" eventid="1087" gender="F" number="3" order="3"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1152" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1153" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1154" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1155" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1156" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1157" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1158" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1159" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1160" agemax="14" agemin="14" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="10:35:00" heatid="1802" number="1" order="1"
                                    status="OFFICIAL" />
                                <HEAT daytime="10:35:00" heatid="1803" number="2" order="2"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
                        </EVENT>
                        <EVENT daytime="10:35:00" eventid="1089" gender="M" number="4" order="4"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1161" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1162" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1163" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1164" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1165" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1166" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1167" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1168" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1169" agemax="14" agemin="14" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="10:35:00" heatid="1804" number="1" order="1"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
                        </EVENT>
                        <EVENT daytime="10:40:00" eventid="1091" gender="F" number="5" order="5"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1170" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1171" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1172" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1173" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1174" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1175" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1176" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1177" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1178" agemax="14" agemin="14" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="10:40:00" heatid="1805" number="1" order="1"
                                    status="OFFICIAL" />
                                <HEAT daytime="10:40:00" heatid="1806" number="2" order="2"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE code="25 СП" distance="25" name="25m На спине" relaycount="1"
                                stroke="UNKNOWN" swimstyleid="103" />
                        </EVENT>
                        <EVENT daytime="10:40:00" eventid="1093" gender="M" number="6" order="6"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1179" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1180" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1181" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1182" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1183" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1184" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1185" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1186" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1187" agemax="14" agemin="14" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="10:40:00" heatid="1807" number="1" order="1"
                                    status="OFFICIAL" />
                                <HEAT daytime="10:45:00" heatid="1808" number="2" order="2"
                                    status="OFFICIAL" />
                                <HEAT daytime="10:45:00" heatid="1809" number="3" order="3"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
                        </EVENT>
                        <EVENT daytime="10:45:00" eventid="1095" gender="F" number="7" order="7"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1188" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1189" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1190" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1191" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1192" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1193" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1194" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1195" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1196" agemax="14" agemin="14" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="10:45:00" heatid="1810" number="1" order="1"
                                    status="OFFICIAL" />
                                <HEAT daytime="10:45:00" heatid="1811" number="2" order="2"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
                        </EVENT>
                        <EVENT daytime="10:50:00" eventid="1099" gender="M" number="8" order="8"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1197" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1198" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1199" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1200" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1201" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1202" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1203" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1204" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1205" agemax="14" agemin="14" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="10:50:00" heatid="1812" number="1" order="1"
                                    status="OFFICIAL" />
                                <HEAT daytime="10:50:00" heatid="1813" number="2" order="2"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
                        </EVENT>
                        <EVENT daytime="10:50:00" eventid="1101" gender="F" number="9" order="9"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1206" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1207" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1208" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1209" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1210" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1211" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1212" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1213" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1214" agemax="14" agemin="14" />
                                <AGEGROUP agegroupid="1762" agemax="15" agemin="15" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="10:50:00" heatid="1814" number="1" order="1"
                                    status="OFFICIAL" />
                                <HEAT daytime="10:55:00" heatid="1815" number="2" order="2"
                                    status="OFFICIAL" />
                                <HEAT daytime="10:55:00" heatid="1816" number="3" order="3"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
                        </EVENT>
                        <EVENT daytime="10:55:00" eventid="1103" gender="M" number="10" order="10"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1215" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1216" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1217" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1218" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1219" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1220" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1221" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1222" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1223" agemax="14" agemin="14" />
                                <AGEGROUP agegroupid="1722" agemax="-1" agemin="15" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="10:55:00" heatid="1817" number="1" order="1"
                                    status="OFFICIAL" />
                                <HEAT daytime="11:00:00" heatid="1818" number="2" order="2"
                                    status="OFFICIAL" />
                                <HEAT daytime="11:00:00" heatid="1819" number="3" order="3"
                                    status="OFFICIAL" />
                                <HEAT daytime="11:05:00" heatid="1820" number="4" order="4"
                                    status="OFFICIAL" />
                                <HEAT daytime="11:05:00" heatid="1821" number="5" order="5"
                                    status="OFFICIAL" />
                                <HEAT daytime="11:05:00" heatid="1822" number="6" order="6"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
                        </EVENT>
                        <EVENT daytime="11:05:00" eventid="1105" gender="F" number="11" order="11"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1224" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1225" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1226" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1227" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1228" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1229" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1230" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1231" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1232" agemax="14" agemin="14" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="11:05:00" heatid="1823" number="1" order="1"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
                        </EVENT>
                        <EVENT daytime="11:10:00" eventid="1107" gender="M" number="12" order="12"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1233" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1234" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1235" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1236" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1237" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1238" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1239" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1240" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1241" agemax="14" agemin="14" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="11:10:00" heatid="1824" number="1" order="1"
                                    status="OFFICIAL" />
                                <HEAT daytime="11:10:00" heatid="1825" number="2" order="2"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
                        </EVENT>
                        <EVENT daytime="11:10:00" eventid="1110" gender="F" number="13" order="13"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1242" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1243" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1244" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1245" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1246" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1247" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1248" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1249" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1250" agemax="14" agemin="14" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="11:10:00" heatid="1826" number="1" order="1"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
                        </EVENT>
                        <EVENT daytime="11:15:00" eventid="1112" gender="M" number="14" order="14"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1251" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1252" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1253" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1254" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1255" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1256" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1257" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1258" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1259" agemax="14" agemin="14" />
                                <AGEGROUP agegroupid="1723" agemax="-1" agemin="15" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="11:15:00" heatid="1827" number="1" order="1"
                                    status="OFFICIAL" />
                                <HEAT daytime="11:15:00" heatid="1828" number="2" order="2"
                                    status="OFFICIAL" />
                                <HEAT daytime="11:20:00" heatid="1829" number="3" order="3"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
                        </EVENT>
                        <EVENT daytime="11:20:00" eventid="1114" gender="F" number="15" order="15"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1260" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1261" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1262" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1263" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1264" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1265" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1266" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1267" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1268" agemax="14" agemin="14" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="11:20:00" heatid="1830" number="1" order="1"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
                        </EVENT>
                        <EVENT daytime="11:20:00" eventid="1116" gender="M" number="16" order="16"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1269" agemax="6" agemin="6" />
                                <AGEGROUP agegroupid="1270" agemax="7" agemin="7" />
                                <AGEGROUP agegroupid="1271" agemax="8" agemin="8" />
                                <AGEGROUP agegroupid="1272" agemax="9" agemin="9" />
                                <AGEGROUP agegroupid="1273" agemax="10" agemin="10" />
                                <AGEGROUP agegroupid="1274" agemax="11" agemin="11" />
                                <AGEGROUP agegroupid="1275" agemax="12" agemin="12" />
                                <AGEGROUP agegroupid="1276" agemax="13" agemin="13" />
                                <AGEGROUP agegroupid="1277" agemax="14" agemin="14" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="11:20:00" heatid="1831" number="1" order="1"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
                        </EVENT>
                    </EVENTS>
                </SESSION>
                <SESSION date="2025-02-02T00:00:00" daytime="11:20:00" number="2">
                    <EVENTS>
                        <EVENT daytime="11:20:00" eventid="1119" gender="F" number="17" order="1"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1120" agemax="-1" agemin="15" />
                            </AGEGROUPS>
                            <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
                        </EVENT>
                        <EVENT daytime="11:20:00" eventid="1121" gender="M" number="18" order="2"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1278" agemax="-1" agemin="15" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="11:20:00" heatid="1832" number="1" order="1"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
                        </EVENT>
                        <EVENT daytime="11:20:00" eventid="1123" gender="F" number="19" order="3"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1279" agemax="-1" agemin="15" />
                            </AGEGROUPS>
                            <SWIMSTYLE code="25 БР" distance="25" name="25m Брасс" relaycount="1"
                                stroke="UNKNOWN" swimstyleid="105" />
                        </EVENT>
                        <EVENT daytime="11:20:00" eventid="1125" gender="M" number="20" order="4"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1280" agemax="-1" agemin="15" />
                            </AGEGROUPS>
                            <SWIMSTYLE code="25 БР" distance="25" name="25m Брасс" relaycount="1"
                                stroke="UNKNOWN" swimstyleid="105" />
                        </EVENT>
                        <EVENT daytime="11:20:00" eventid="1127" gender="F" number="21" order="5"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1281" agemax="-1" agemin="15" />
                            </AGEGROUPS>
                            <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
                        </EVENT>
                        <EVENT daytime="11:20:00" eventid="1129" gender="M" number="22" order="6"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1282" agemax="-1" agemin="15" />
                            </AGEGROUPS>
                            <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
                        </EVENT>
                        <EVENT daytime="11:20:00" eventid="1131" gender="F" number="23" order="7"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1283" agemax="-1" agemin="15" />
                            </AGEGROUPS>
                            <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
                        </EVENT>
                        <EVENT daytime="11:20:00" eventid="1133" gender="M" number="24" order="8"
                            preveventid="-1" round="TIM">
                            <AGEGROUPS>
                                <AGEGROUP agegroupid="1284" agemax="-1" agemin="15" />
                            </AGEGROUPS>
                            <HEATS>
                                <HEAT daytime="11:20:00" heatid="1833" number="1" order="1"
                                    status="OFFICIAL" />
                            </HEATS>
                            <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
                        </EVENT>
                    </EVENTS>
                </SESSION>
            </SESSIONS>
        </MEET>
    </MEETS>
</LENEX>